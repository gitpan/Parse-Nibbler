

module 

	hello   

	(
                portname,  otherport
		,yetanotherport



			);


input     portname;

output
	otherport;

inout	yetanotherport;

 	modulename instance_name_1 ( port1[7:0], {port2a, port2b, port2c}, port3[12], , ,  port4 );

			endmodule





