
module my_mod (port1, port2, port3);

input port1;
output port3;

my_mod inst_name ( .port1({connector1,signal2}), .port2(1'b1) );

endmodule



