
module my_mod 
(
port1, port2, port3
)

;


input port1;

output port2;
inout port3;

my_mod inst_name ( );

endmodule



